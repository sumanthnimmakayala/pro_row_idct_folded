// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
/*
 *-------------------------------------------------------------
 *
 * user_proj_example
 *
 * This is an example of a (trivially simple) user project,
 * showing how the user project can connect to the logic
 * analyzer, the wishbone bus, and the I/O pads.
 *
 * This project generates an integer count, which is output
 * on the user area GPIO pads (digital output only).  The
 * wishbone connection allows the project to be controlled
 * (start and stop) from the management SoC program.
 *
 * See the testbenches in directory "mprj_counter" for the
 * example programs that drive this user project.  The three
 * testbenches are "io_ports", "la_test1", and "la_test2".
 *
 *-------------------------------------------------------------
 */

module user_proj_example #(
    parameter BITS = 32
)(
`ifdef USE_POWER_PINS
    inout vccd1,	// User area 1 1.8V supply
    inout vssd1,	// User area 1 digital ground
`endif

    // Wishbone Slave ports (WB MI A)
    input wb_clk_i,
    input wb_rst_i,
    input wbs_stb_i,
    input wbs_cyc_i,
    input wbs_we_i,
    input [3:0] wbs_sel_i,
    input [31:0] wbs_dat_i,
    input [31:0] wbs_adr_i,
    output wbs_ack_o,
    output [31:0] wbs_dat_o,

    // Logic Analyzer Signals
    input  [127:0] la_data_in,
    output [127:0] la_data_out,
    input  [127:0] la_oenb,

    // IOs
    input  [`MPRJ_IO_PADS-1:0] io_in,
    output [`MPRJ_IO_PADS-1:0] io_out,
    output [`MPRJ_IO_PADS-1:0] io_oeb,

    // IRQ
    output [2:0] irq
);
    wire clk;
    wire rst;

    wire [`MPRJ_IO_PADS-1:0] io_in;
    wire [`MPRJ_IO_PADS-1:0] io_out;
    wire [`MPRJ_IO_PADS-1:0] io_oeb;

    wire [31:0] rdata; 
    wire [31:0] wdata;
    wire [BITS-1:0] count;

    wire valid;
    wire [3:0] wstrb;
    wire [31:0] la_write;

    // WB MI A
    assign valid = wbs_cyc_i && wbs_stb_i; 
    assign wstrb = wbs_sel_i & {4{wbs_we_i}};
    assign wbs_dat_o = rdata;
    assign wdata = wbs_dat_i;

    // IO
    assign io_out = count;
    assign io_oeb = {(`MPRJ_IO_PADS-1){rst}};

    // IRQ
    assign irq = 3'b000;	// Unused

    // LA
    assign la_data_out = {{(127-BITS){1'b0}}, count};
    // Assuming LA probes [63:32] are for controlling the count register  
    assign la_write = ~la_oenb[63:32] & ~{BITS{valid}};
    // Assuming LA probes [65:64] are for controlling the count clk & reset  
    assign clk = (~la_oenb[64]) ? la_data_in[64]: wb_clk_i;
    assign rst = (~la_oenb[65]) ? la_data_in[65]: wb_rst_i;

pro_row_idct_folded dut(

i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
s,se,

ou20s,ou21s,ou22s,ou23s,ou24s,ou25s,ou26s,ou27s,ou28s,ou29s,ou210s,ou211s,ou212s,ou213s,ou214s,ou215s,
ou20,ou21,ou22,ou23,ou24,ou25,ou26,ou27,ou28,ou29,ou210,ou211,ou212,ou213,ou214,ou215,

ou40s,ou41s,ou42s,ou43s,ou44s,ou45s,ou46s,ou47s,
ou40,ou41,ou42,ou43,ou44,ou45,ou46,ou47,

ou80s,ou81s,ou82s,ou83s,
ou80,ou81,ou82,ou83,

ou160s,ou161s,
ou160,ou161,

ou320s,
ou320

);

endmodule

//proposed 32-point configurable IntegerDCT for row process in folded architecture

//`include "block_complete_row_folded.v"
//`include "cell_sign.v"
//`include "adder40.v"

module pro_row_idct_folded(

i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
s,se,

ou20s,ou21s,ou22s,ou23s,ou24s,ou25s,ou26s,ou27s,ou28s,ou29s,ou210s,ou211s,ou212s,ou213s,ou214s,ou215s,
ou20,ou21,ou22,ou23,ou24,ou25,ou26,ou27,ou28,ou29,ou210,ou211,ou212,ou213,ou214,ou215,

ou40s,ou41s,ou42s,ou43s,ou44s,ou45s,ou46s,ou47s,
ou40,ou41,ou42,ou43,ou44,ou45,ou46,ou47,

ou80s,ou81s,ou82s,ou83s,
ou80,ou81,ou82,ou83,

ou160s,ou161s,
ou160,ou161,

ou320s,
ou320

);

output ou20s,ou21s,ou22s,ou23s,ou24s,ou25s,ou26s,ou27s,ou28s,ou29s,ou210s,ou211s,ou212s,ou213s,ou214s,ou215s,
ou40s,ou41s,ou42s,ou43s,ou44s,ou45s,ou46s,ou47s,
ou80s,ou81s,ou82s,ou83s,
ou160s,ou161s,
ou320s;

output [39:0] ou20,ou21,ou22,ou23,ou24,ou25,ou26,ou27,ou28,ou29,ou210,ou211,ou212,ou213,ou214,ou215,
ou40,ou41,ou42,ou43,ou44,ou45,ou46,ou47,
ou80,ou81,ou82,ou83,
ou160,ou161,
ou320;

input i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s;
input [39:0] i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31;

input [4:0] s;
input [2:0] se;

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

wire [39:0] o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,o10,o11,o12,o13,o14,o15,o16,o17,o18,o19,o20,o21,o22,o23,o24,o25,o26,o27,o28,o29,o30,o31;
wire o0s,o1s,o2s,o3s,o4s,o5s,o6s,o7s,o8s,o9s,o10s,o11s,o12s,o13s,o14s,o15s,o16s,o17s,o18s,o19s,o20s,o21s,o22s,o23s,o24s,o25s,o26s,o27s,o28s,o29s,o30s,o31s;

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp0(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o0

);

cell_sign cc0(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o0s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp1(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o1

);

cell_sign cc1(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o1s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp2(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o2

);

cell_sign cc2(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o2s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp3(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o3

);

cell_sign cc3(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o3s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp4(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o4

);

cell_sign cc4(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o4s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp5(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o5

);

cell_sign cc5(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o5s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp6(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o6

);

cell_sign cc6(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o6s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp7(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o7

);

cell_sign cc7(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o7s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp8(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o8

);

cell_sign cc8(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o8s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp9(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o9

);

cell_sign cc9(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o9s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp10(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o10

);

cell_sign cc10(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o10s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp11(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o11

);

cell_sign cc11(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o11s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp12(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o12

);

cell_sign cc12(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o12s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp13(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o13

);

cell_sign cc13(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o13s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp14(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o14

);

cell_sign cc14(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o14s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp15(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o15

);

cell_sign cc15(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o15s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp16(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o16

);

cell_sign cc16(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o16s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp17(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o17

);

cell_sign cc17(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o17s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp18(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o18

);

cell_sign cc18(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o18s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp19(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o19

);

cell_sign cc19(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o19s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp20(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o20

);

cell_sign cc20(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o20s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp21(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o21

);

cell_sign cc21(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o21s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp22(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o22

);

cell_sign cc22(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o22s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp23(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o23

);

cell_sign cc23(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o23s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp24(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o24

);

cell_sign cc24(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o24s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp25(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o25

);

cell_sign cc25(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o25s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp26(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o26

);

cell_sign cc26(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o26s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp27(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o27

);

cell_sign cc27(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o27s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp28(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o28

);

cell_sign cc28(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o28s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp29(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o29

);

cell_sign cc29(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o29s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp30(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o30

);

cell_sign cc30(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o30s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_folded pp31(

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,
i0,i1,i2,i3,i4,i5,i6,i7,
i0,i1,i2,i3,
i0,i1,

s,se,o31

);

cell_sign cc31(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o31s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

wire ou20s,ou21s,ou22s,ou23s,ou24s,ou25s,ou26s,ou27s,ou28s,ou29s,ou210s,ou211s,ou212s,ou213s,ou214s,ou215s,
ou40s,ou41s,ou42s,ou43s,ou44s,ou45s,ou46s,ou47s,
ou80s,ou81s,ou82s,ou83s,
ou160s,ou161s,
ou320s;

wire [39:0] ou20,ou21,ou22,ou23,ou24,ou25,ou26,ou27,ou28,ou29,ou210,ou211,ou212,ou213,ou214,ou215,
ou40,ou41,ou42,ou43,ou44,ou45,ou46,ou47,
ou80,ou81,ou82,ou83,
ou160,ou161,
ou320;

//first level of tree of adders

adder40 ad10(o0s,o0,o1s,o1,ou20s,ou20);
adder40 ad11(o2s,o2,o3s,o3,ou21s,ou21);
adder40 ad12(o4s,o4,o5s,o5,ou22s,ou22);
adder40 ad13(o6s,o6,o7s,o7,ou23s,ou23);
adder40 ad14(o8s,o8,o9s,o9,ou24s,ou24);
adder40 ad15(o10s,o10,o11s,o11,ou25s,ou25);
adder40 ad16(o12s,o12,o13s,o13,ou26s,ou26);
adder40 ad17(o14s,o14,o15s,o15,ou27s,ou27);
adder40 ad18(o16s,o16,o17s,o17,ou28s,ou28);
adder40 ad19(o18s,o18,o19s,o19,ou29s,ou29);
adder40 ad110(o20s,o20,o21s,o21,ou210s,ou210);
adder40 ad111(o22s,o22,o23s,o23,ou211s,ou211);
adder40 ad112(o24s,o24,o25s,o25,ou212s,ou212);
adder40 ad113(o26s,o26,o27s,o27,ou213s,ou213);
adder40 ad114(o28s,o28,o29s,o29,ou214s,ou214);
adder40 ad115(o30s,o30,o31s,o31,ou215s,ou215);

//second level of tree of adders

adder40 ad20(ou20s,ou20,ou21s,ou21,ou40s,ou40);
adder40 ad21(ou22s,ou22,ou23s,ou23,ou41s,ou41);
adder40 ad22(ou24s,ou24,ou25s,ou25,ou42s,ou42);
adder40 ad23(ou26s,ou26,ou27s,ou27,ou43s,ou43);
adder40 ad24(ou28s,ou28,ou29s,ou29,ou44s,ou44);
adder40 ad25(ou210s,ou210,ou211s,ou211,ou45s,ou45);
adder40 ad26(ou212s,ou212,ou213s,ou213,ou46s,ou46);
adder40 ad27(ou214s,ou214,ou215s,ou215,ou47s,ou47);

//third level of tree of adders

adder40 ad30(ou40s,ou40,ou41s,ou41,ou80s,ou80);
adder40 ad31(ou42s,ou42,ou43s,ou43,ou81s,ou81);
adder40 ad32(ou44s,ou44,ou45s,ou45,ou82s,ou82);
adder40 ad33(ou46s,ou46,ou47s,ou47,ou83s,ou83);

//fourth level of tree of adders

adder40 ad40(ou80s,ou80,ou81s,ou81,ou160s,ou160);
adder40 ad41(ou82s,ou82,ou83s,ou83,ou161s,ou161);

//fifth level of tree of adders

adder40 ad50(ou160s,ou160,ou161s,ou161,ou320s,ou320);

endmodule


//40 bit fixed point adder

//`include "recurse40.v"
//`include "kgp.v"
//`include "kgp_carry.v"
//`include "recursive_stage1.v"

module adder40(as,a,bs,in_b,rrs,rr);

input as,bs;
input [39:0] a,in_b;
output rrs;
output [39:0] rr;

reg rrs;
reg [39:0] rr;
wire z;
assign z=as^bs;
wire cout,cout1;

wire [39:0] r1,b1,b2;
assign b1=(~in_b);

recurse40 c0(b2,cout1,b1,40'd1);

reg [39:0] b;

always@(z or in_b or b2)
	begin
		if(z==0)
			b=in_b;
		else if (z==1)
			b=b2;
	end
	
recurse40 c1(r1,cout,a,b);

wire cout2;
wire [39:0] r11,r22;
assign r11=(~r1);
recurse40 c2(r22,cout2,r11,40'd1);

reg carry;
always@(r1 or cout or z or as or bs or r22)
 begin
	if(z==0)	
		begin
			rrs=as;
			rr=r1;
			carry=cout;
		end
	else if (z==1 && cout==1)
		begin	
			rrs=as;
			rr=r1;
			carry=1'b0;
		end
	else if (z==1 && cout==0)
		begin
			rrs=(~as);
			rr=r22;
			carry=1'b0;
		end
 end

endmodule


/*`include "mux32to1_1.v"
`include "mux16to1_1.v"
`include "mux8to1_1.v"
`include "mux4to1_1.v"
`include "mux2to1_1.v"
`include "mux5to1_1.v"*/

//cell used for sign in Integer DCT 

module cell_sign(i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,s,se,out);

input i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31;
input [4:0] s;
input [2:0] se;
output out;

wire out1,out2,out3,out4,out5;

wire si0,si1,si2,si3,si4,si5,si6,si7,si8,si9,si10,si11,si12,si13,si14,si15,si16,si17,si18,si19,si20,si21,si22,si23,si24,si25,si26,si27,si28,si29,si30,si31;

assign si0=i0^1'b0;
assign si1=i1^1'b0;
assign si2=i2^1'b0;
assign si3=i3^1'b0;
assign si4=i4^1'b0;
assign si5=i5^1'b0;
assign si6=i6^1'b0;
assign si7=i7^1'b0;
assign si8=i8^1'b0;
assign si9=i9^1'b0;
assign si10=i10^1'b0;
assign si11=i11^1'b0;
assign si12=i12^1'b0;
assign si13=i13^1'b0;
assign si14=i14^1'b0;
assign si15=i15^1'b0;
assign si16=i16^1'b0;
assign si17=i17^1'b0;
assign si18=i18^1'b0;
assign si19=i19^1'b0;
assign si20=i20^1'b0;
assign si21=i21^1'b0;
assign si22=i22^1'b0;
assign si23=i23^1'b0;
assign si24=i24^1'b0;
assign si25=i25^1'b0;
assign si26=i26^1'b0;
assign si27=i27^1'b0;
assign si28=i28^1'b0;
assign si29=i29^1'b0;
assign si30=i30^1'b0;
assign si31=i31^1'b0;

mux32to1_1 mu1(out1,si0,si1,si2,si3,si4,si5,si6,si7,si8,si9,si10,si11,si12,si13,si14,si15,si16,si17,si18,si19,si20,si21,si22,si23,si24,si25,si26,si27,si28,si29,si30,si31,s[4],s[3],s[2],s[1],s[0]);
mux16to1_1 mu2(out2,si0,si1,si2,si3,si4,si5,si6,si7,si8,si9,si10,si11,si12,si13,si14,si15,s[3:0]);
mux8to1_1 mmu3(out3,si0,si1,si2,si3,si4,si5,si6,si7,s[2:0]);
mux4to1_1 mmu4(out4,si0,si1,si2,si3,s[1:0]);
mux2to1_1 mmu5(out5,si0,si1,s[0]);
mux5to1_1 mmu6(out,out1,out2,out3,out4,out5,se);

endmodule


//The complete block used for row process in parallel architecture

//`include "cell_row_folded.v"
//`include "block_row_folded.v"

module block_complete_row_folded(

i00,i01,i02,i03,i04,i05,i06,i07,i08,i09,i010,i011,i012,i013,i014,i015,i016,i017,i018,i019,i020,i021,i022,i023,i024,i025,i026,i027,i028,i029,i030,i031,
n00,n01,n02,n03,n04,n05,n06,n07,n08,n09,n010,n011,n012,n013,n014,n015,
m00,m01,m02,m03,m04,m05,m06,m07,
o00,o01,o02,o03,
p00,p01,

i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i110,i111,i112,i113,i114,i115,i116,i117,i118,i119,i120,i121,i122,i123,i124,i125,i126,i127,i128,i129,i130,i131,
n10,n11,n12,n13,n14,n15,n16,n17,n18,n19,n110,n111,n112,n113,n114,n115,
m10,m11,m12,m13,m14,m15,m16,m17,
o10,o11,o12,o13,
p10,p11,

i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i210,i211,i212,i213,i214,i215,i216,i217,i218,i219,i220,i221,i222,i223,i224,i225,i226,i227,i228,i229,i230,i231,
n20,n21,n22,n23,n24,n25,n26,n27,n28,n29,n210,n211,n212,n213,n214,n215,
m20,m21,m22,m23,m24,m25,m26,m27,
o20,o21,o22,o23,
p20,p21,

i30,i31,i32,i33,i34,i35,i36,i37,i38,i39,i310,i311,i312,i313,i314,i315,i316,i317,i318,i319,i320,i321,i322,i323,i324,i325,i326,i327,i328,i329,i330,i331,
n30,n31,n32,n33,n34,n35,n36,n37,n38,n39,n310,n311,n312,n313,n314,n315,
m30,m31,m32,m33,m34,m35,m36,m37,
o30,o31,o32,o33,
p30,p31,

i40,i41,i42,i43,i44,i45,i46,i47,i48,i49,i410,i411,i412,i413,i414,i415,i416,i417,i418,i419,i420,i421,i422,i423,i424,i425,i426,i427,i428,i429,i430,i431,
n40,n41,n42,n43,n44,n45,n46,n47,n48,n49,n410,n411,n412,n413,n414,n415,
m40,m41,m42,m43,m44,m45,m46,m47,
o40,o41,o42,o43,
p40,p41,

s,se,out

);

output [39:0] out;

input [4:0] s;
input [2:0] se;

input [39:0] i00,i01,i02,i03,i04,i05,i06,i07,i08,i09,i010,i011,i012,i013,i014,i015,i016,i017,i018,i019,i020,i021,i022,i023,i024,i025,i026,i027,i028,i029,i030,i031,
n00,n01,n02,n03,n04,n05,n06,n07,n08,n09,n010,n011,n012,n013,n014,n015,
m00,m01,m02,m03,m04,m05,m06,m07,
o00,o01,o02,o03,
p00,p01,

i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i110,i111,i112,i113,i114,i115,i116,i117,i118,i119,i120,i121,i122,i123,i124,i125,i126,i127,i128,i129,i130,i131,
n10,n11,n12,n13,n14,n15,n16,n17,n18,n19,n110,n111,n112,n113,n114,n115,
m10,m11,m12,m13,m14,m15,m16,m17,
o10,o11,o12,o13,
p10,p11,

i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i210,i211,i212,i213,i214,i215,i216,i217,i218,i219,i220,i221,i222,i223,i224,i225,i226,i227,i228,i229,i230,i231,
n20,n21,n22,n23,n24,n25,n26,n27,n28,n29,n210,n211,n212,n213,n214,n215,
m20,m21,m22,m23,m24,m25,m26,m27,
o20,o21,o22,o23,
p20,p21,

i30,i31,i32,i33,i34,i35,i36,i37,i38,i39,i310,i311,i312,i313,i314,i315,i316,i317,i318,i319,i320,i321,i322,i323,i324,i325,i326,i327,i328,i329,i330,i331,
n30,n31,n32,n33,n34,n35,n36,n37,n38,n39,n310,n311,n312,n313,n314,n315,
m30,m31,m32,m33,m34,m35,m36,m37,
o30,o31,o32,o33,
p30,p31,

i40,i41,i42,i43,i44,i45,i46,i47,i48,i49,i410,i411,i412,i413,i414,i415,i416,i417,i418,i419,i420,i421,i422,i423,i424,i425,i426,i427,i428,i429,i430,i431,
n40,n41,n42,n43,n44,n45,n46,n47,n48,n49,n410,n411,n412,n413,n414,n415,
m40,m41,m42,m43,m44,m45,m46,m47,
o40,o41,o42,o43,
p40,p41;

wire [39:0] b0,b1,b2,b3,b4;

cell_row_folded c0(i00,i01,i02,i03,i04,i05,i06,i07,i08,i09,i010,i011,i012,i013,i014,i015,i016,i017,i018,i019,i020,i021,i022,i023,i024,i025,i026,i027,i028,i029,i030,i031,
n00,n01,n02,n03,n04,n05,n06,n07,n08,n09,n010,n011,n012,n013,n014,n015,
m00,m01,m02,m03,m04,m05,m06,m07,
o00,o01,o02,o03,
p00,p01,
s,se,b0

);

cell_row_folded c1(i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i110,i111,i112,i113,i114,i115,i116,i117,i118,i119,i120,i121,i122,i123,i124,i125,i126,i127,i128,i129,i130,i131,
n10,n11,n12,n13,n14,n15,n16,n17,n18,n19,n110,n111,n112,n113,n114,n115,
m10,m11,m12,m13,m14,m15,m16,m17,
o10,o11,o12,o13,
p10,p11,
s,se,b1

);

cell_row_folded c2(i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i210,i211,i212,i213,i214,i215,i216,i217,i218,i219,i220,i221,i222,i223,i224,i225,i226,i227,i228,i229,i230,i231,
n20,n21,n22,n23,n24,n25,n26,n27,n28,n29,n210,n211,n212,n213,n214,n215,
m20,m21,m22,m23,m24,m25,m26,m27,
o20,o21,o22,o23,
p20,p21,
s,se,b2

);

cell_row_folded c3(i30,i31,i32,i33,i34,i35,i36,i37,i38,i39,i310,i311,i312,i313,i314,i315,i316,i317,i318,i319,i320,i321,i322,i323,i324,i325,i326,i327,i328,i329,i330,i331,
n30,n31,n32,n33,n34,n35,n36,n37,n38,n39,n310,n311,n312,n313,n314,n315,
m30,m31,m32,m33,m34,m35,m36,m37,
o30,o31,o32,o33,
p30,p31,
s,se,b3

);

cell_row_folded c4(i40,i41,i42,i43,i44,i45,i46,i47,i48,i49,i410,i411,i412,i413,i414,i415,i416,i417,i418,i419,i420,i421,i422,i423,i424,i425,i426,i427,i428,i429,i430,i431,
n40,n41,n42,n43,n44,n45,n46,n47,n48,n49,n410,n411,n412,n413,n414,n415,
m40,m41,m42,m43,m44,m45,m46,m47,
o40,o41,o42,o43,
p40,p41,
s,se,b4

);

block_row_folded block(b0,b1,b2,b3,b4,out);

endmodule

/*`include "mux32to1_40.v"
`include "mux16to1_40.v"
`include "mux8to1_40.v"
`include "mux4to1_40.v"
`include "mux2to1_40.v"
`include "mux5to1_40.v"*/

//cell used for row process in folded architecture of Integer DCT

module cell_row_folded(i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
n0,n1,n2,n3,n4,n5,n6,n7,n8,n9,n10,n11,n12,n13,n14,n15,
m0,m1,m2,m3,m4,m5,m6,m7,
o0,o1,o2,o3,
p0,p1,
s,se,out

);

input [39:0] i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
n0,n1,n2,n3,n4,n5,n6,n7,n8,n9,n10,n11,n12,n13,n14,n15,
m0,m1,m2,m3,m4,m5,m6,m7,
o0,o1,o2,o3,
p0,p1;

input [4:0] s;
input [2:0] se;
output [39:0] out;

wire [39:0] out1,out2,out3,out4,out5;

mux32to1_40 mu1(out1,i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,s[4],s[3],s[2],s[1],s[0]);
mux16to1_40 mu2(out2,n0,n1,n2,n3,n4,n5,n6,n7,n8,n9,n10,n11,n12,n13,n14,n15,s[3:0]);
mux8to1_40 mmu3(out3,m0,m1,m2,m3,m4,m5,m6,m7,s[2:0]);
mux4to1_40 mmu4(out4,o0,o1,o2,o3,s[1:0]);
mux2to1_40 mmu5(out5,p0,p1,s[0]);
mux5to1_40 mmu6(out,out1,out2,out3,out4,out5,se);

endmodule


/*
`include "halfadd.v"
`include "fulladd.v"
`include "kgp.v"
`include "kgp_carry.v"
`include "recursive_stage1.v"
`include "recurse40.v"*/

//block used for row process in parallel architecture

module block_row_folded(i0,i1,i2,i3,i4,out);

input [39:0] i0,i1,i2,i3,i4;
output [39:0] out;

wire [39:0] sum1h,sum11h,sum2h;
wire carry1h,carry11h,carry2h,carry;

recurse40 rr1(sum1h,carry1h,i0,i1);
recurse40 rr2(sum11h,carry11h,i2,i3);
recurse40 rr3(sum2h,carry2h,sum1h,sum11h); 
recurse40 rr4(out,carry,sum2h,i4); 

endmodule


module kgp(a,b,y);

input a,b;
output [1:0] y;
//reg [1:0] y;

//always@(a or b)
//begin
//case({a,b})
//2'b00:y=2'b00;  //kill
//2'b11:y=2'b11;	  //generate
//2'b01:y=2'b01;	//propagate
//2'b10:y=2'b01;  //propagate
//endcase   //y[1]=ab  y[0]=a+b  
//end

assign y[0]=a | b;
assign y[1]=a & b;

endmodule




module kgp_carry(a,b,carry);

input [1:0] a,b;
output carry;
reg carry;

always@(a or b)
begin
case(a)
2'b00:carry=1'b0;  
2'b11:carry=1'b1;
2'b01:carry=b[0];
2'b10:carry=b[0];
default:carry=1'bx;
endcase
end

/*wire carry;

wire f,g;
assign g=a[0] & a[1];
assign f=a[0] ^ a[1];

assign carry=g|(b[0] & f);*/

endmodule


module recursive_stage1(a,b,y);

input [1:0] a,b;
output [1:0] y;

wire [1:0] y;
wire b0;
not n1(b0,b[1]);
wire f,g0,g1;
and a1(f,b[0],b[1]);
and a2(g0,b0,b[0],a[0]);
and a3(g1,b0,b[0],a[1]);

or o1(y[0],f,g0);
or o2(y[1],f,g1);

//reg [1:0] y;
//always@(a or b)
//begin
//case(b)
//2'b00:y=2'b00;  
//2'b11:y=2'b11;
//2'b01:y=a;
//default:y=2'bx;
//endcase
//end

//always@(a or b)
//begin
//if(b==2'b00)
//	y=2'b00;  
//else if (b==2'b11)
//	y=2'b11;
//else if (b==2'b01)
//	y=a;
//end

//wire x;
//assign x=a[0] ^ b[0];
//always@(a or b or x)
//begin
//case(x)
//1'b0:y[0]=b[0];  
//1'b1:y[0]=a[0]; 
//endcase
//end
//
//always@(a or b or x)
//begin
//case(x)
//1'b0:y[1]=b[1];  
//1'b1:y[1]=a[1];
//endcase
//end


//always@(a or b)
//begin
//if (b==2'b00)
//	y=2'b00; 
//else if (b==2'b11)	
//	y=2'b11;
//else if (b==2'b01 && a==2'b00)
//	y=2'b00;
//else if (b==2'b01 && a==2'b11)
//	y=2'b11;
//else if (b==2'b01 && a==2'b01)
//	y=2'b01;
//end

endmodule

//40 bit recursive doubling technique

module recurse40(sum,carry,a,b); 

output [39:0] sum;
output  carry;
input [39:0] a,b;

wire [81:0] x;

assign x[1:0]=2'b00;  // kgp generation

kgp a00(a[0],b[0],x[3:2]);
kgp a01(a[1],b[1],x[5:4]);
kgp a02(a[2],b[2],x[7:6]);
kgp a03(a[3],b[3],x[9:8]);
kgp a04(a[4],b[4],x[11:10]);
kgp a05(a[5],b[5],x[13:12]);
kgp a06(a[6],b[6],x[15:14]);
kgp a07(a[7],b[7],x[17:16]);
kgp a08(a[8],b[8],x[19:18]);
kgp a09(a[9],b[9],x[21:20]);
kgp a10(a[10],b[10],x[23:22]);
kgp a11(a[11],b[11],x[25:24]);
kgp a12(a[12],b[12],x[27:26]);
kgp a13(a[13],b[13],x[29:28]);
kgp a14(a[14],b[14],x[31:30]);
kgp a15(a[15],b[15],x[33:32]);
kgp a16(a[16],b[16],x[35:34]);
kgp a17(a[17],b[17],x[37:36]);
kgp a18(a[18],b[18],x[39:38]);
kgp a19(a[19],b[19],x[41:40]);
kgp a20(a[20],b[20],x[43:42]);
kgp a21(a[21],b[21],x[45:44]);
kgp a22(a[22],b[22],x[47:46]);
kgp a23(a[23],b[23],x[49:48]);
kgp a24(a[24],b[24],x[51:50]);
kgp a25(a[25],b[25],x[53:52]);
kgp a26(a[26],b[26],x[55:54]);
kgp a27(a[27],b[27],x[57:56]);
kgp a28(a[28],b[28],x[59:58]);
kgp a29(a[29],b[29],x[61:60]);
kgp a30(a[30],b[30],x[63:62]);
kgp a31(a[31],b[31],x[65:64]);
kgp a32(a[32],b[32],x[67:66]);
kgp a33(a[33],b[33],x[69:68]);
kgp a34(a[34],b[34],x[71:70]);
kgp a35(a[35],b[35],x[73:72]);
kgp a36(a[36],b[36],x[75:74]);
kgp a37(a[37],b[37],x[77:76]);
kgp a38(a[38],b[38],x[79:78]);
kgp a39(a[39],b[39],x[81:80]);

wire [79:0] x1;  //recursive doubling stage 1
assign x1[1:0]=x[1:0];

recursive_stage1 s00(x[1:0],x[3:2],x1[3:2]);
recursive_stage1 s01(x[3:2],x[5:4],x1[5:4]);
recursive_stage1 s02(x[5:4],x[7:6],x1[7:6]);
recursive_stage1 s03(x[7:6],x[9:8],x1[9:8]);
recursive_stage1 s04(x[9:8],x[11:10],x1[11:10]);
recursive_stage1 s05(x[11:10],x[13:12],x1[13:12]);
recursive_stage1 s06(x[13:12],x[15:14],x1[15:14]);
recursive_stage1 s07(x[15:14],x[17:16],x1[17:16]);
recursive_stage1 s08(x[17:16],x[19:18],x1[19:18]);
recursive_stage1 s09(x[19:18],x[21:20],x1[21:20]);
recursive_stage1 s10(x[21:20],x[23:22],x1[23:22]);
recursive_stage1 s11(x[23:22],x[25:24],x1[25:24]);
recursive_stage1 s12(x[25:24],x[27:26],x1[27:26]);
recursive_stage1 s13(x[27:26],x[29:28],x1[29:28]);
recursive_stage1 s14(x[29:28],x[31:30],x1[31:30]);
recursive_stage1 s15(x[31:30],x[33:32],x1[33:32]);
recursive_stage1 s16(x[33:32],x[35:34],x1[35:34]);
recursive_stage1 s17(x[35:34],x[37:36],x1[37:36]);
recursive_stage1 s18(x[37:36],x[39:38],x1[39:38]);
recursive_stage1 s19(x[39:38],x[41:40],x1[41:40]);
recursive_stage1 s20(x[41:40],x[43:42],x1[43:42]);
recursive_stage1 s21(x[43:42],x[45:44],x1[45:44]);
recursive_stage1 s22(x[45:44],x[47:46],x1[47:46]);
recursive_stage1 s23(x[47:46],x[49:48],x1[49:48]);
recursive_stage1 s24(x[49:48],x[51:50],x1[51:50]);
recursive_stage1 s25(x[51:50],x[53:52],x1[53:52]);
recursive_stage1 s26(x[53:52],x[55:54],x1[55:54]);
recursive_stage1 s27(x[55:54],x[57:56],x1[57:56]);
recursive_stage1 s28(x[57:56],x[59:58],x1[59:58]);
recursive_stage1 s29(x[59:58],x[61:60],x1[61:60]);
recursive_stage1 s30(x[61:60],x[63:62],x1[63:62]);
recursive_stage1 s31(x[63:62],x[65:64],x1[65:64]);
recursive_stage1 s32(x[65:64],x[67:66],x1[67:66]);
recursive_stage1 s33(x[67:66],x[69:68],x1[69:68]);
recursive_stage1 s34(x[69:68],x[71:70],x1[71:70]);
recursive_stage1 s35(x[71:70],x[73:72],x1[73:72]);
recursive_stage1 s36(x[73:72],x[75:74],x1[75:74]);
recursive_stage1 s37(x[75:74],x[77:76],x1[77:76]);
recursive_stage1 s38(x[77:76],x[79:78],x1[79:78]);

wire [79:0] x2;  //recursive doubling stage2
assign x2[3:0]=x1[3:0];

recursive_stage1 s101(x1[1:0],x1[5:4],x2[5:4]);
recursive_stage1 s102(x1[3:2],x1[7:6],x2[7:6]);
recursive_stage1 s103(x1[5:4],x1[9:8],x2[9:8]);
recursive_stage1 s104(x1[7:6],x1[11:10],x2[11:10]);
recursive_stage1 s105(x1[9:8],x1[13:12],x2[13:12]);
recursive_stage1 s106(x1[11:10],x1[15:14],x2[15:14]);
recursive_stage1 s107(x1[13:12],x1[17:16],x2[17:16]);
recursive_stage1 s108(x1[15:14],x1[19:18],x2[19:18]);
recursive_stage1 s109(x1[17:16],x1[21:20],x2[21:20]);
recursive_stage1 s110(x1[19:18],x1[23:22],x2[23:22]);
recursive_stage1 s111(x1[21:20],x1[25:24],x2[25:24]);
recursive_stage1 s112(x1[23:22],x1[27:26],x2[27:26]);
recursive_stage1 s113(x1[25:24],x1[29:28],x2[29:28]);
recursive_stage1 s114(x1[27:26],x1[31:30],x2[31:30]);
recursive_stage1 s115(x1[29:28],x1[33:32],x2[33:32]);
recursive_stage1 s116(x1[31:30],x1[35:34],x2[35:34]);
recursive_stage1 s117(x1[33:32],x1[37:36],x2[37:36]);
recursive_stage1 s118(x1[35:34],x1[39:38],x2[39:38]);
recursive_stage1 s119(x1[37:36],x1[41:40],x2[41:40]);
recursive_stage1 s120(x1[39:38],x1[43:42],x2[43:42]);
recursive_stage1 s121(x1[41:40],x1[45:44],x2[45:44]);
recursive_stage1 s122(x1[43:42],x1[47:46],x2[47:46]);
recursive_stage1 s123(x1[45:44],x1[49:48],x2[49:48]);
recursive_stage1 s124(x1[47:46],x1[51:50],x2[51:50]);
recursive_stage1 s125(x1[49:48],x1[53:52],x2[53:52]);
recursive_stage1 s126(x1[51:50],x1[55:54],x2[55:54]);
recursive_stage1 s127(x1[53:52],x1[57:56],x2[57:56]);
recursive_stage1 s128(x1[55:54],x1[59:58],x2[59:58]);
recursive_stage1 s129(x1[57:56],x1[61:60],x2[61:60]);
recursive_stage1 s130(x1[59:58],x1[63:62],x2[63:62]);
recursive_stage1 s131(x1[61:60],x1[65:64],x2[65:64]);
recursive_stage1 s132(x1[63:62],x1[67:66],x2[67:66]);
recursive_stage1 s133(x1[65:64],x1[69:68],x2[69:68]);
recursive_stage1 s134(x1[67:66],x1[71:70],x2[71:70]);
recursive_stage1 s135(x1[69:68],x1[73:72],x2[73:72]);
recursive_stage1 s136(x1[71:70],x1[75:74],x2[75:74]);
recursive_stage1 s137(x1[73:72],x1[77:76],x2[77:76]);
recursive_stage1 s138(x1[75:74],x1[79:78],x2[79:78]);

wire [79:0] x3;  //recursive doubling stage3
assign x3[7:0]=x2[7:0];

recursive_stage1 s203(x2[1:0],x2[9:8],x3[9:8]);
recursive_stage1 s204(x2[3:2],x2[11:10],x3[11:10]);
recursive_stage1 s205(x2[5:4],x2[13:12],x3[13:12]);
recursive_stage1 s206(x2[7:6],x2[15:14],x3[15:14]);
recursive_stage1 s207(x2[9:8],x2[17:16],x3[17:16]);
recursive_stage1 s208(x2[11:10],x2[19:18],x3[19:18]);
recursive_stage1 s209(x2[13:12],x2[21:20],x3[21:20]);
recursive_stage1 s210(x2[15:14],x2[23:22],x3[23:22]);
recursive_stage1 s211(x2[17:16],x2[25:24],x3[25:24]);
recursive_stage1 s212(x2[19:18],x2[27:26],x3[27:26]);
recursive_stage1 s213(x2[21:20],x2[29:28],x3[29:28]);
recursive_stage1 s214(x2[23:22],x2[31:30],x3[31:30]);
recursive_stage1 s215(x2[25:24],x2[33:32],x3[33:32]);
recursive_stage1 s216(x2[27:26],x2[35:34],x3[35:34]);
recursive_stage1 s217(x2[29:28],x2[37:36],x3[37:36]);
recursive_stage1 s218(x2[31:30],x2[39:38],x3[39:38]);
recursive_stage1 s219(x2[33:32],x2[41:40],x3[41:40]);
recursive_stage1 s220(x2[35:34],x2[43:42],x3[43:42]);
recursive_stage1 s221(x2[37:36],x2[45:44],x3[45:44]);
recursive_stage1 s222(x2[39:38],x2[47:46],x3[47:46]);
recursive_stage1 s223(x2[41:40],x2[49:48],x3[49:48]);
recursive_stage1 s224(x2[43:42],x2[51:50],x3[51:50]);
recursive_stage1 s225(x2[45:44],x2[53:52],x3[53:52]);
recursive_stage1 s226(x2[47:46],x2[55:54],x3[55:54]);
recursive_stage1 s227(x2[49:48],x2[57:56],x3[57:56]);
recursive_stage1 s228(x2[51:50],x2[59:58],x3[59:58]);
recursive_stage1 s229(x2[53:52],x2[61:60],x3[61:60]);
recursive_stage1 s230(x2[55:54],x2[63:62],x3[63:62]);
recursive_stage1 s231(x2[57:56],x2[65:64],x3[65:64]);
recursive_stage1 s232(x2[59:58],x2[67:66],x3[67:66]);
recursive_stage1 s233(x2[61:60],x2[69:68],x3[69:68]);
recursive_stage1 s234(x2[63:62],x2[71:70],x3[71:70]);
recursive_stage1 s235(x2[65:64],x2[73:72],x3[73:72]);
recursive_stage1 s236(x2[67:66],x2[75:74],x3[75:74]);
recursive_stage1 s237(x2[69:68],x2[77:76],x3[77:76]);
recursive_stage1 s238(x2[71:70],x2[79:78],x3[79:78]);

wire [79:0] x4;  //recursive doubling stage 4
assign x4[15:0]=x3[15:0];

recursive_stage1 s307(x3[1:0],x3[17:16],x4[17:16]);
recursive_stage1 s308(x3[3:2],x3[19:18],x4[19:18]);
recursive_stage1 s309(x3[5:4],x3[21:20],x4[21:20]);
recursive_stage1 s310(x3[7:6],x3[23:22],x4[23:22]);
recursive_stage1 s311(x3[9:8],x3[25:24],x4[25:24]);
recursive_stage1 s312(x3[11:10],x3[27:26],x4[27:26]);
recursive_stage1 s313(x3[13:12],x3[29:28],x4[29:28]);
recursive_stage1 s314(x3[15:14],x3[31:30],x4[31:30]);
recursive_stage1 s315(x3[17:16],x3[33:32],x4[33:32]);
recursive_stage1 s316(x3[19:18],x3[35:34],x4[35:34]);
recursive_stage1 s317(x3[21:20],x3[37:36],x4[37:36]);
recursive_stage1 s318(x3[23:22],x3[39:38],x4[39:38]);
recursive_stage1 s319(x3[25:24],x3[41:40],x4[41:40]);
recursive_stage1 s320(x3[27:26],x3[43:42],x4[43:42]);
recursive_stage1 s321(x3[29:28],x3[45:44],x4[45:44]);
recursive_stage1 s322(x3[31:30],x3[47:46],x4[47:46]);
recursive_stage1 s323(x3[33:32],x3[49:48],x4[49:48]);
recursive_stage1 s324(x3[35:34],x3[51:50],x4[51:50]);
recursive_stage1 s325(x3[37:36],x3[53:52],x4[53:52]);
recursive_stage1 s326(x3[39:38],x3[55:54],x4[55:54]);
recursive_stage1 s327(x3[41:40],x3[57:56],x4[57:56]);
recursive_stage1 s328(x3[43:42],x3[59:58],x4[59:58]);
recursive_stage1 s329(x3[45:44],x3[61:60],x4[61:60]);
recursive_stage1 s330(x3[47:46],x3[63:62],x4[63:62]);
recursive_stage1 s331(x3[49:48],x3[65:64],x4[65:64]);
recursive_stage1 s332(x3[51:50],x3[67:66],x4[67:66]);
recursive_stage1 s333(x3[53:52],x3[69:68],x4[69:68]);
recursive_stage1 s334(x3[55:54],x3[71:70],x4[71:70]);
recursive_stage1 s335(x3[57:56],x3[73:72],x4[73:72]);
recursive_stage1 s336(x3[59:58],x3[75:74],x4[75:74]);
recursive_stage1 s337(x3[61:60],x3[77:76],x4[77:76]);
recursive_stage1 s338(x3[63:62],x3[79:78],x4[79:78]);

wire [79:0] x5;  //recursive doubling stage 5
assign x5[31:0]=x4[31:0];

recursive_stage1 s415(x4[1:0],x4[33:32],x5[33:32]);
recursive_stage1 s416(x4[3:2],x4[35:34],x5[35:34]);
recursive_stage1 s417(x4[5:4],x4[37:36],x5[37:36]);
recursive_stage1 s418(x4[7:6],x4[39:38],x5[39:38]);
recursive_stage1 s419(x4[9:8],x4[41:40],x5[41:40]);
recursive_stage1 s420(x4[11:10],x4[43:42],x5[43:42]);
recursive_stage1 s421(x4[13:12],x4[45:44],x5[45:44]);
recursive_stage1 s422(x4[15:14],x4[47:46],x5[47:46]);
recursive_stage1 s423(x4[17:16],x4[49:48],x5[49:48]);
recursive_stage1 s424(x4[19:18],x4[51:50],x5[51:50]);
recursive_stage1 s425(x4[21:20],x4[53:52],x5[53:52]);
recursive_stage1 s426(x4[23:22],x4[55:54],x5[55:54]);
recursive_stage1 s427(x4[25:24],x4[57:56],x5[57:56]);
recursive_stage1 s428(x4[27:26],x4[59:58],x5[59:58]);
recursive_stage1 s429(x4[29:28],x4[61:60],x5[61:60]);
recursive_stage1 s430(x4[31:30],x4[63:62],x5[63:62]);
recursive_stage1 s431(x4[33:32],x4[65:64],x5[65:64]);
recursive_stage1 s432(x4[35:34],x4[67:66],x5[67:66]);
recursive_stage1 s433(x4[37:36],x4[69:68],x5[69:68]);
recursive_stage1 s434(x4[39:38],x4[71:70],x5[71:70]);
recursive_stage1 s435(x4[41:40],x4[73:72],x5[73:72]);
recursive_stage1 s436(x4[43:42],x4[75:74],x5[75:74]);
recursive_stage1 s437(x4[45:44],x4[77:76],x5[77:76]);
recursive_stage1 s438(x4[47:46],x4[79:78],x5[79:78]);

wire [79:0] x6;  // recursive doubling stage 6
assign x6[63:0]=x5[63:0];

recursive_stage1 s531(x5[1:0],x5[65:64],x6[65:64]);
recursive_stage1 s532(x5[3:2],x5[67:66],x6[67:66]);
recursive_stage1 s533(x5[5:4],x5[69:68],x6[69:68]);
recursive_stage1 s534(x5[7:6],x5[71:70],x6[71:70]);
recursive_stage1 s535(x5[9:8],x5[73:72],x6[73:72]);
recursive_stage1 s536(x5[11:10],x5[75:74],x6[75:74]);
recursive_stage1 s537(x5[13:12],x5[77:76],x6[77:76]);
recursive_stage1 s538(x5[15:14],x5[79:78],x6[79:78]);

// final sum and carry

assign sum[0]=a[0]^b[0]^x6[0];
assign sum[1]=a[1]^b[1]^x6[2];
assign sum[2]=a[2]^b[2]^x6[4];
assign sum[3]=a[3]^b[3]^x6[6];
assign sum[4]=a[4]^b[4]^x6[8];
assign sum[5]=a[5]^b[5]^x6[10];
assign sum[6]=a[6]^b[6]^x6[12];
assign sum[7]=a[7]^b[7]^x6[14];
assign sum[8]=a[8]^b[8]^x6[16];
assign sum[9]=a[9]^b[9]^x6[18];
assign sum[10]=a[10]^b[10]^x6[20];
assign sum[11]=a[11]^b[11]^x6[22];
assign sum[12]=a[12]^b[12]^x6[24];
assign sum[13]=a[13]^b[13]^x6[26];
assign sum[14]=a[14]^b[14]^x6[28];
assign sum[15]=a[15]^b[15]^x6[30];
assign sum[16]=a[16]^b[16]^x6[32];
assign sum[17]=a[17]^b[17]^x6[34];
assign sum[18]=a[18]^b[18]^x6[36];
assign sum[19]=a[19]^b[19]^x6[38];
assign sum[20]=a[20]^b[20]^x6[40];
assign sum[21]=a[21]^b[21]^x6[42];
assign sum[22]=a[22]^b[22]^x6[44];
assign sum[23]=a[23]^b[23]^x6[46];
assign sum[24]=a[24]^b[24]^x6[48];
assign sum[25]=a[25]^b[25]^x6[50];
assign sum[26]=a[26]^b[26]^x6[52];
assign sum[27]=a[27]^b[27]^x6[54];
assign sum[28]=a[28]^b[28]^x6[56];
assign sum[29]=a[29]^b[29]^x6[58];
assign sum[30]=a[30]^b[30]^x6[60];
assign sum[31]=a[31]^b[31]^x6[62];
assign sum[32]=a[32]^b[32]^x6[64];
assign sum[33]=a[33]^b[33]^x6[66];
assign sum[34]=a[34]^b[34]^x6[68];
assign sum[35]=a[35]^b[35]^x6[70];
assign sum[36]=a[36]^b[36]^x6[72];
assign sum[37]=a[37]^b[37]^x6[74];
assign sum[38]=a[38]^b[38]^x6[76];
assign sum[39]=a[39]^b[39]^x6[79];

kgp_carry kkc(x[81:80],x6[79:78],carry);

endmodule


//mux32to1

module mux32to1_40(out,i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,s4,s3,s2,s1,s0);
input [39:0] i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31;
input s4,s3,s2,s1,s0;
output [39:0] out;

//level 1 

reg [39:0] out;

always@(i0 or i1 or i2 or i3 or i4 or i5 or i6 or i7 or i8 or i9 or i10 or i11 or i12 or i13 or i14 or i15 or i16 or i17 or i18 or i19 or i20 or i21 or i22 or i23 or i24 or i25 or i26 or i27 or i28 or i29 or i30 or i31 or s4 or s3 or s2 or s1 or s0)
begin 
case({s4,s3,s2,s1,s0})
5'b00000: out = i0;
5'b00001: out = i1;
5'b00010: out = i2;
5'b00011: out = i3;
5'b00100: out = i4;
5'b00101: out = i5;
5'b00110: out = i6;
5'b00111: out = i7;
5'b01000: out = i8;
5'b01001: out = i9;
5'b01010: out = i10;
5'b01011: out = i11;
5'b01100: out = i12;
5'b01101: out = i13;
5'b01110: out = i14;
5'b01111: out = i15;
5'b10000: out = i16;
5'b10001: out = i17;
5'b10010: out = i18;
5'b10011: out = i19;
5'b10100: out = i20;
5'b10101: out = i21;
5'b10110: out = i22;
5'b10111: out = i23;
5'b11000: out = i24;
5'b11001: out = i25;
5'b11010: out = i26;
5'b11011: out = i27;
5'b11100: out = i28;
5'b11101: out = i29;
5'b11110: out = i30;
5'b11111: out = i31;
default: out = 40'bx;
endcase
end 


endmodule

//mux16to1

module mux16to1_40(o,i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,s);

input [39:0] i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15;
input [3:0] s;
output [39:0] o;
reg [39:0] o;

always@(i0 or i1 or i2 or i3 or i4 or i5 or i6 or i7 or i8 or i9 or i10 or i11 or i12 or i13 or i14 or i15 or s)
	begin
		case(s)
		 4'b0000:o=i0;
		 4'b0001:o=i1;
		 4'b0010:o=i2;
		 4'b0011:o=i3;
		 4'b0100:o=i4;
		 4'b0101:o=i5;
		 4'b0110:o=i6;
		 4'b0111:o=i7;
		 4'b1000:o=i8;
		 4'b1001:o=i9;
		 4'b1010:o=i10;
		 4'b1011:o=i11;
		 4'b1100:o=i12;
		 4'b1101:o=i13;
		 4'b1110:o=i14;
		 4'b1111:o=i15;
		 //default:o=1'bx;
		endcase
	end


endmodule



//mux8to1

module mux8to1_40(o,i0,i1,i2,i3,i4,i5,i6,i7,s);

input [39:0] i0,i1,i2,i3,i4,i5,i6,i7;
input [2:0] s;
output [39:0] o;
reg [39:0] o;

always@(i0 or i1 or i2 or i3 or i4 or i5 or i6 or i7 or s)
	begin
		case(s)
		 3'b000:o=i0;
		 3'b001:o=i1;
		 3'b010:o=i2;
		 3'b011:o=i3;
		 3'b100:o=i4;
		 3'b101:o=i5;
		 3'b110:o=i6;
		 3'b111:o=i7;
		 //default:o=1'bx;
		endcase
	end


endmodule


//mux4to1

module mux4to1_40(y,in0,in1,in2,in3,sel);

input [39:0] in0,in1,in2,in3;
input [1:0] sel;
output [39:0] y;

reg [39:0] y;
always@(in0 or in1 or in2 or in3 or sel)
begin
case(sel)
2'b00:y=in0;  
2'b01:y=in1;
2'b10:y=in2;	
2'b11:y=in3;  
//default:y=1'bx;
endcase   
end


endmodule



//2-to-1 multiplexer design

module mux2to1_40(out,i1,i2,s);

input [39:0] i1,i2;
input s;
output [39:0] out;
reg [39:0] out;

always@(i1 or i2 or s)
	begin
	 case(s)
	  1'b0:out=i1;
	  1'b1:out=i2;
	 endcase
	end

endmodule


//mux5 to 1

module mux5to1_40(o,o1,o2,o3,o4,o5,dir);

input [2:0] dir;
input [39:0] o1,o2,o3,o4,o5;
output [39:0] o;

reg [39:0] o;

always@(o1 or o2 or o3 or o4 or o5 or dir)
	begin
	 case(dir)
	  3'b000: o=o1;
	  3'b001: o=o2;
	  3'b010: o=o3;
	  3'b011: o=o4;
	  3'b100: o=o5;	  
	default: o = 1'bx;
	 endcase
	end

endmodule



//mux32to1

module mux32to1_1(out,i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,s4,s3,s2,s1,s0);
input i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,s4,s3,s2,s1,s0;
output out;

//level 1 

reg out;

always@(i0 or i1 or i2 or i3 or i4 or i5 or i6 or i7 or i8 or i9 or i10 or i11 or i12 or i13 or i14 or i15 or i16 or i17 or i18 or i19 or i20 or i21 or i22 or i23 or i24 or i25 or i26 or i27 or i28 or i29 or i30 or i31 or s4 or s3 or s2 or s1 or s0)
begin 
case({s4,s3,s2,s1,s0})
5'b00000: out = i0;
5'b00001: out = i1;
5'b00010: out = i2;
5'b00011: out = i3;
5'b00100: out = i4;
5'b00101: out = i5;
5'b00110: out = i6;
5'b00111: out = i7;
5'b01000: out = i8;
5'b01001: out = i9;
5'b01010: out = i10;
5'b01011: out = i11;
5'b01100: out = i12;
5'b01101: out = i13;
5'b01110: out = i14;
5'b01111: out = i15;
5'b10000: out = i16;
5'b10001: out = i17;
5'b10010: out = i18;
5'b10011: out = i19;
5'b10100: out = i20;
5'b10101: out = i21;
5'b10110: out = i22;
5'b10111: out = i23;
5'b11000: out = i24;
5'b11001: out = i25;
5'b11010: out = i26;
5'b11011: out = i27;
5'b11100: out = i28;
5'b11101: out = i29;
5'b11110: out = i30;
5'b11111: out = i31;
default: out = 1'bx;
endcase
end 


endmodule


//mux16to1

module mux16to1_1(o,i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,s);

input i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15;
input [3:0] s;
output o;
reg o;

always@(i0 or i1 or i2 or i3 or i4 or i5 or i6 or i7 or i8 or i9 or i10 or i11 or i12 or i13 or i14 or i15 or s)
	begin
		case(s)
		 4'b0000:o=i0;
		 4'b0001:o=i1;
		 4'b0010:o=i2;
		 4'b0011:o=i3;
		 4'b0100:o=i4;
		 4'b0101:o=i5;
		 4'b0110:o=i6;
		 4'b0111:o=i7;
		 4'b1000:o=i8;
		 4'b1001:o=i9;
		 4'b1010:o=i10;
		 4'b1011:o=i11;
		 4'b1100:o=i12;
		 4'b1101:o=i13;
		 4'b1110:o=i14;
		 4'b1111:o=i15;
		 //default:o=1'bx;
		endcase
	end


endmodule



//mux8to1

module mux8to1_1(o,i0,i1,i2,i3,i4,i5,i6,i7,s);

input i0,i1,i2,i3,i4,i5,i6,i7;
input [2:0] s;
output o;
reg o;

always@(i0 or i1 or i2 or i3 or i4 or i5 or i6 or i7 or s)
	begin
		case(s)
		 3'b000:o=i0;
		 3'b001:o=i1;
		 3'b010:o=i2;
		 3'b011:o=i3;
		 3'b100:o=i4;
		 3'b101:o=i5;
		 3'b110:o=i6;
		 3'b111:o=i7;
		 //default:o=1'bx;
		endcase
	end


endmodule


//mux4to1

module mux4to1_1(y,in0,in1,in2,in3,sel);

input in0,in1,in2,in3;
input [1:0] sel;
output y;

reg y;
always@(in0 or in1 or in2 or in3 or sel)
begin
case(sel)
2'b00:y=in0;  
2'b01:y=in1;
2'b10:y=in2;	
2'b11:y=in3;  
//default:y=1'bx;
endcase   
end

endmodule


//2 to 1 multiplexer design

module mux2to1_1(out,i1,i2,s);

input i1,i2,s;
output out;
reg out;

always@(i1 or i2 or s)
	begin
	 case(s)
	  1'b0:out=i1;
	  1'b1:out=i2;
	 endcase
	end

endmodule



//mux5 to 1

module mux5to1_1(o,o1,o2,o3,o4,o5,dir);

input [2:0] dir;
input o1,o2,o3,o4,o5;
output o;

reg o;

always@(o1 or o2 or o3 or o4 or o5 or dir)
	begin
	 case(dir)
	  3'b000: o=o1;
	  3'b001: o=o2;
	  3'b010: o=o3;
	  3'b011: o=o4;
	  3'b100: o=o5;
	  
	default: o = 1'bx;
	 endcase
	end

endmodule

//32-point proposed Integer DCT using folded architecture 

//`include "folded_buffer_pro.v"
//`include "pro_row_idct_folded.v"

module idct_proposed_folded(

i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
s,se,ss,clk,reset,
se0,se1,se2,se3,se4,se5,se6,se7,se8,se9,se10,se11,se12,se13,se14,se15,se16,se17,se18,se19,se20,se21,se22,se23,se24,se25,se26,se27,se28,se29,se30,se31,

oo0,oo1,oo2,oo3,oo4,oo5,oo6,oo7,oo8,oo9,oo10,oo11,oo12,oo13,oo14,oo15,oo16,oo17,oo18,oo19,oo20,oo21,oo22,oo23,oo24,oo25,oo26,oo27,oo28,oo29,oo30,oo31,
oo0s,oo1s,oo2s,oo3s,oo4s,oo5s,oo6s,oo7s,oo8s,oo9s,oo10s,oo11s,oo12s,oo13s,oo14s,oo15s,oo16s,oo17s,oo18s,oo19s,oo20s,oo21s,oo22s,oo23s,
oo24s,oo25s,oo26s,oo27s,oo28s,oo29s,oo30s,oo31s


);

input clk,reset;

input i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s;
input [7:0] i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31;

input [4:0] s;
input [2:0] se;
input ss;//ss=0 for row process and ss=1 for column process

input se0,se1,se2,se3,se4,se5,se6,se7,se8,se9,se10,se11,se12,se13,se14,se15,se16,se17,se18,se19,se20,se21,se22,se23,se24,se25,se26,se27,se28,se29,se30,se31;

output [39:0] oo0,oo1,oo2,oo3,oo4,oo5,oo6,oo7,oo8,oo9,oo10,oo11,oo12,oo13,oo14,oo15,oo16,oo17,oo18,oo19,oo20,oo21,oo22,oo23,oo24,oo25,oo26,oo27,oo28,oo29,oo30,oo31;
output oo0s,oo1s,oo2s,oo3s,oo4s,oo5s,oo6s,oo7s,oo8s,oo9s,oo10s,oo11s,oo12s,oo13s,oo14s,oo15s,oo16s,oo17s,oo18s,oo19s,oo20s,oo21s,oo22s,
oo23s,oo24s,oo25s,oo26s,oo27s,oo28s,oo29s,oo30s,oo31s;

//selection of row and column processes

wire in0s,in1s,in2s,in3s,in4s,in5s,in6s,in7s,in8s,in9s,in10s,in11s,in12s,in13s,in14s,in15s,in16s,in17s,in18s,in19s,in20s,in21s,in22s,in23s,in24s,in25s,in26s,in27s,in28s,in29s,in30s,in31s;
wire [39:0] in0,in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31;

mux2to1_41 mu0({in0s,in0},{i0s,32'd0,i0},{oo0s,oo0},ss);
mux2to1_41 mu1({in1s,in1},{i1s,32'd0,i1},{oo1s,oo1},ss);
mux2to1_41 mu2({in2s,in2},{i2s,32'd0,i2},{oo2s,oo2},ss);
mux2to1_41 mu3({in3s,in3},{i3s,32'd0,i3},{oo3s,oo3},ss);
mux2to1_41 mu4({in4s,in4},{i4s,32'd0,i4},{oo4s,oo4},ss);
mux2to1_41 mu5({in5s,in5},{i5s,32'd0,i5},{oo5s,oo5},ss);
mux2to1_41 mu6({in6s,in6},{i6s,32'd0,i6},{oo6s,oo6},ss);
mux2to1_41 mu7({in7s,in7},{i7s,32'd0,i7},{oo7s,oo7},ss);
mux2to1_41 mu8({in8s,in8},{i8s,32'd0,i8},{oo8s,oo8},ss);
mux2to1_41 mu9({in9s,in9},{i9s,32'd0,i9},{oo9s,oo9},ss);
mux2to1_41 mu10({in10s,in10},{i10s,32'd0,i10},{oo10s,oo10},ss);
mux2to1_41 mu11({in11s,in11},{i11s,32'd0,i11},{oo11s,oo11},ss);
mux2to1_41 mu12({in12s,in12},{i12s,32'd0,i12},{oo12s,oo12},ss);
mux2to1_41 mu13({in13s,in13},{i13s,32'd0,i13},{oo13s,oo13},ss);
mux2to1_41 mu14({in14s,in14},{i14s,32'd0,i14},{oo14s,oo14},ss);
mux2to1_41 mu15({in15s,in15},{i15s,32'd0,i15},{oo15s,oo15},ss);
mux2to1_41 mu16({in16s,in16},{i16s,32'd0,i16},{oo16s,oo16},ss);
mux2to1_41 mu17({in17s,in17},{i17s,32'd0,i17},{oo17s,oo17},ss);
mux2to1_41 mu18({in18s,in18},{i18s,32'd0,i18},{oo18s,oo18},ss);
mux2to1_41 mu19({in19s,in19},{i19s,32'd0,i19},{oo19s,oo19},ss);
mux2to1_41 mu20({in20s,in20},{i20s,32'd0,i20},{oo20s,oo20},ss);
mux2to1_41 mu21({in21s,in21},{i21s,32'd0,i21},{oo21s,oo21},ss);
mux2to1_41 mu22({in22s,in22},{i22s,32'd0,i22},{oo22s,oo22},ss);
mux2to1_41 mu23({in23s,in23},{i23s,32'd0,i23},{oo23s,oo23},ss);
mux2to1_41 mu24({in24s,in24},{i24s,32'd0,i24},{oo24s,oo24},ss);
mux2to1_41 mu25({in25s,in25},{i25s,32'd0,i25},{oo25s,oo25},ss);
mux2to1_41 mu26({in26s,in26},{i26s,32'd0,i26},{oo26s,oo26},ss);
mux2to1_41 mu27({in27s,in27},{i27s,32'd0,i27},{oo27s,oo27},ss);
mux2to1_41 mu28({in28s,in28},{i28s,32'd0,i28},{oo28s,oo28},ss);
mux2to1_41 mu29({in29s,in29},{i29s,32'd0,i29},{oo29s,oo29},ss);
mux2to1_41 mu30({in30s,in30},{i30s,32'd0,i30},{oo30s,oo30},ss);
mux2to1_41 mu31({in31s,in31},{i31s,32'd0,i31},{oo31s,oo31},ss);

//row and column process

wire ou20s,ou21s,ou22s,ou23s,ou24s,ou25s,ou26s,ou27s,ou28s,ou29s,ou210s,ou211s,ou212s,ou213s,ou214s,ou215s,
ou40s,ou41s,ou42s,ou43s,ou44s,ou45s,ou46s,ou47s,
ou80s,ou81s,ou82s,ou83s,
ou160s,ou161s,
ou320s;

wire [39:0] ou20,ou21,ou22,ou23,ou24,ou25,ou26,ou27,ou28,ou29,ou210,ou211,ou212,ou213,ou214,ou215,
ou40,ou41,ou42,ou43,ou44,ou45,ou46,ou47,
ou80,ou81,ou82,ou83,
ou160,ou161,
ou320;

pro_row_idct_folded mod_1(

in0s,in1s,in2s,in3s,in4s,in5s,in6s,in7s,in8s,in9s,in10s,in11s,in12s,in13s,in14s,in15s,in16s,in17s,in18s,in19s,in20s,in21s,in22s,in23s,in24s,in25s,in26s,in27s,in28s,in29s,in30s,in31s,
in0,in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,
s,se,

ou20s,ou21s,ou22s,ou23s,ou24s,ou25s,ou26s,ou27s,ou28s,ou29s,ou210s,ou211s,ou212s,ou213s,ou214s,ou215s,
ou20,ou21,ou22,ou23,ou24,ou25,ou26,ou27,ou28,ou29,ou210,ou211,ou212,ou213,ou214,ou215,

ou40s,ou41s,ou42s,ou43s,ou44s,ou45s,ou46s,ou47s,
ou40,ou41,ou42,ou43,ou44,ou45,ou46,ou47,

ou80s,ou81s,ou82s,ou83s,
ou80,ou81,ou82,ou83,

ou160s,ou161s,
ou160,ou161,

ou320s,
ou320

);

//transpose buffer

wire out20s,out21s,out22s,out23s,out24s,out25s,out26s,out27s,out28s,out29s,out210s,out211s,out212s,out213s,out214s,out215s,
out40s,out41s,out42s,out43s,out44s,out45s,out46s,out47s,
out80s,out81s,out82s,out83s,
out160s,out161s,
out320s;

wire [39:0] out20,out21,out22,out23,out24,out25,out26,out27,out28,out29,out210,out211,out212,out213,out214,out215,
out40,out41,out42,out43,out44,out45,out46,out47,
out80,out81,out82,out83,
out160,out161,
out320;

assign {out20s,out20}={ou20s,16'd0,ou20};
assign {out21s,out21}={ou21s,16'd0,ou21};
assign {out22s,out22}={ou22s,16'd0,ou22};
assign {out23s,out23}={ou23s,16'd0,ou23};
assign {out24s,out24}={ou24s,16'd0,ou24};
assign {out25s,out25}={ou25s,16'd0,ou25};
assign {out26s,out26}={ou26s,16'd0,ou26};
assign {out27s,out27}={ou27s,16'd0,ou27};
assign {out28s,out28}={ou28s,16'd0,ou28};
assign {out29s,out29}={ou29s,16'd0,ou29};
assign {out210s,out210}={ou210s,16'd0,ou210};
assign {out211s,out211}={ou211s,16'd0,ou211};
assign {out212s,out212}={ou212s,16'd0,ou212};
assign {out213s,out213}={ou213s,16'd0,ou213};
assign {out214s,out214}={ou214s,16'd0,ou214};
assign {out215s,out215}={ou215s,16'd0,ou215};
assign {out40s,out40}={ou40s,16'd0,ou40};
assign {out41s,out41}={ou41s,16'd0,ou41};
assign {out42s,out42}={ou42s,16'd0,ou42};
assign {out43s,out43}={ou43s,16'd0,ou43};
assign {out44s,out44}={ou44s,16'd0,ou44};
assign {out45s,out45}={ou45s,16'd0,ou45};
assign {out46s,out46}={ou46s,16'd0,ou46};
assign {out47s,out47}={ou47s,16'd0,ou47};
assign {out80s,out80}={ou80s,16'd0,ou80};
assign {out81s,out81}={ou81s,16'd0,ou81};
assign {out82s,out82}={ou82s,16'd0,ou82};
assign {out83s,out83}={ou83s,16'd0,ou83};
assign {out160s,out160}={ou160s,16'd0,ou160};
assign {out161s,out161}={ou161s,16'd0,ou161};
assign {out320s,out320}={ou320s,16'd0,ou320};

folded_buffer_pro mod_2(

out20s,out21s,out22s,out23s,out24s,out25s,out26s,out27s,out28s,out29s,out210s,out211s,out212s,out213s,out214s,out215s,
out20,out21,out22,out23,out24,out25,out26,out27,out28,out29,out210,out211,out212,out213,out214,out215,

out40s,out41s,out42s,out43s,out44s,out45s,out46s,out47s,
out40,out41,out42,out43,out44,out45,out46,out47,

out80s,out81s,out82s,out83s,
out80,out81,out82,out83,

out160s,out161s,
out160,out161,

out320s,
out320,

se,clk,reset,

se0,se1,se2,se3,se4,se5,se6,se7,se8,se9,se10,se11,se12,se13,se14,se15,se16,se17,se18,se19,se20,se21,se22,se23,se24,se25,se26,se27,se28,se29,se30,se31,

oo0s,oo1s,oo2s,oo3s,oo4s,oo5s,oo6s,oo7s,oo8s,oo9s,oo10s,oo11s,oo12s,oo13s,oo14s,oo15s,oo16s,oo17s,oo18s,oo19s,oo20s,oo21s,oo22s,oo23s,
oo24s,oo25s,oo26s,oo27s,oo28s,oo29s,oo30s,oo31s,
oo0,oo1,oo2,oo3,oo4,oo5,oo6,oo7,oo8,oo9,oo10,oo11,oo12,oo13,oo14,oo15,oo16,oo17,oo18,oo19,oo20,oo21,oo22,oo23,oo24,oo25,oo26,oo27,oo28,oo29,oo30,oo31



);

endmodule


//32x32 buffer with column of multiplexers in proposed Interger DCT parallel architecture

//`include "col_mux_inp_buf_folded_pro.v"
//`include "storage32_41.v"
//`include "mux5_41.v"

module folded_buffer_pro(

ou20s,ou21s,ou22s,ou23s,ou24s,ou25s,ou26s,ou27s,ou28s,ou29s,ou210s,ou211s,ou212s,ou213s,ou214s,ou215s,
ou20,ou21,ou22,ou23,ou24,ou25,ou26,ou27,ou28,ou29,ou210,ou211,ou212,ou213,ou214,ou215,

ou40s,ou41s,ou42s,ou43s,ou44s,ou45s,ou46s,ou47s,
ou40,ou41,ou42,ou43,ou44,ou45,ou46,ou47,

ou80s,ou81s,ou82s,ou83s,
ou80,ou81,ou82,ou83,

ou160s,ou161s,
ou160,ou161,

ou320s,
ou320,

se,clk,reset,

se0,se1,se2,se3,se4,se5,se6,se7,se8,se9,se10,se11,se12,se13,se14,se15,se16,se17,se18,se19,se20,se21,se22,se23,se24,se25,se26,se27,se28,se29,se30,se31,

oo0s,oo1s,oo2s,oo3s,oo4s,oo5s,oo6s,oo7s,oo8s,oo9s,oo10s,oo11s,oo12s,oo13s,oo14s,oo15s,oo16s,oo17s,oo18s,oo19s,oo20s,oo21s,oo22s,oo23s,oo24s,oo25s,oo26s,oo27s,oo28s,oo29s,oo30s,oo31s,
oo0,oo1,oo2,oo3,oo4,oo5,oo6,oo7,oo8,oo9,oo10,oo11,oo12,oo13,oo14,oo15,oo16,oo17,oo18,oo19,oo20,oo21,oo22,oo23,oo24,oo25,oo26,oo27,oo28,oo29,oo30,oo31

);

input clk,reset;

output [39:0] oo0,oo1,oo2,oo3,oo4,oo5,oo6,oo7,oo8,oo9,oo10,oo11,oo12,oo13,oo14,oo15,oo16,oo17,oo18,oo19,oo20,oo21,oo22,oo23,oo24,oo25,oo26,oo27,oo28,oo29,oo30,oo31;
output oo0s,oo1s,oo2s,oo3s,oo4s,oo5s,oo6s,oo7s,oo8s,oo9s,oo10s,oo11s,oo12s,oo13s,oo14s,oo15s,oo16s,oo17s,oo18s,oo19s,oo20s,oo21s,oo22s,oo23s,oo24s,oo25s,oo26s,oo27s,oo28s,oo29s,oo30s,oo31s;

input se0,se1,se2,se3,se4,se5,se6,se7,se8,se9,se10,se11,se12,se13,se14,se15,se16,se17,se18,se19,se20,se21,se22,se23,se24,se25,se26,se27,se28,se29,se30,se31;

input ou20s,ou21s,ou22s,ou23s,ou24s,ou25s,ou26s,ou27s,ou28s,ou29s,ou210s,ou211s,ou212s,ou213s,ou214s,ou215s,
ou40s,ou41s,ou42s,ou43s,ou44s,ou45s,ou46s,ou47s,
ou80s,ou81s,ou82s,ou83s,
ou160s,ou161s,
ou320s;

input [39:0] ou20,ou21,ou22,ou23,ou24,ou25,ou26,ou27,ou28,ou29,ou210,ou211,ou212,ou213,ou214,ou215,
ou40,ou41,ou42,ou43,ou44,ou45,ou46,ou47,
ou80,ou81,ou82,ou83,
ou160,ou161,
ou320;

input [2:0] se;

wire [39:0] o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,o10,o11,o12,o13,o14,o15,o16,o17,o18,o19,o20,o21,o22,o23,o24,o25,o26,o27,o28,o29,o30,o31;
wire o0s,o1s,o2s,o3s,o4s,o5s,o6s,o7s,o8s,o9s,o10s,o11s,o12s,o13s,o14s,o15s,o16s,o17s,o18s,o19s,o20s,o21s,o22s,o23s,o24s,o25s,o26s,o27s,o28s,o29s,o30s,o31s;

col_mux_inp_buf_folded_pro mod1(

ou20s,ou21s,ou22s,ou23s,ou24s,ou25s,ou26s,ou27s,ou28s,ou29s,ou210s,ou211s,ou212s,ou213s,ou214s,ou215s,
ou40s,ou41s,ou42s,ou43s,ou44s,ou45s,ou46s,ou47s,
ou80s,ou81s,ou82s,ou83s,
ou160s,ou161s,
ou320s,

ou20,ou21,ou22,ou23,ou24,ou25,ou26,ou27,ou28,ou29,ou210,ou211,ou212,ou213,ou214,ou215,
ou40,ou41,ou42,ou43,ou44,ou45,ou46,ou47,
ou80,ou81,ou82,ou83,
ou160,ou161,
ou320,

se,

o0s,o1s,o2s,o3s,o4s,o5s,o6s,o7s,o8s,o9s,o10s,o11s,o12s,o13s,o14s,o15s,o16s,o17s,o18s,o19s,o20s,o21s,o22s,o23s,o24s,o25s,o26s,o27s,o28s,o29s,o30s,o31s,
o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,o10,o11,o12,o13,o14,o15,o16,o17,o18,o19,o20,o21,o22,o23,o24,o25,o26,o27,o28,o29,o30,o31

);

wire [40:0] d002,d004,d008,d0016,d0032;
wire [40:0] d012,d014,d018,d0116,d0132;
wire [40:0] d022,d024,d028,d0216,d0232;
wire [40:0] d032,d034,d038,d0316,d0332;
wire [40:0] d042,d044,d048,d0416,d0432;
wire [40:0] d052,d054,d058,d0516,d0532;
wire [40:0] d062,d064,d068,d0616,d0632;
wire [40:0] d072,d074,d078,d0716,d0732;
wire [40:0] d082,d084,d088,d0816,d0832;
wire [40:0] d092,d094,d098,d0916,d0932;


wire [40:0] d102,d104,d108,d1016,d1032;
wire [40:0] d112,d114,d118,d1116,d1132;
wire [40:0] d122,d124,d128,d1216,d1232;
wire [40:0] d132,d134,d138,d1316,d1332;
wire [40:0] d142,d144,d148,d1416,d1432;
wire [40:0] d152,d154,d158,d1516,d1532;
wire [40:0] d162,d164,d168,d1616,d1632;
wire [40:0] d172,d174,d178,d1716,d1732;
wire [40:0] d182,d184,d188,d1816,d1832;
wire [40:0] d192,d194,d198,d1916,d1932;
wire [40:0] d202,d204,d208,d2016,d2032;
wire [40:0] d212,d214,d218,d2116,d2132;
wire [40:0] d222,d224,d228,d2216,d2232;
wire [40:0] d232,d234,d238,d2316,d2332;
wire [40:0] d242,d244,d248,d2416,d2432;
wire [40:0] d252,d254,d258,d2516,d2532;
wire [40:0] d262,d264,d268,d2616,d2632;
wire [40:0] d272,d274,d278,d2716,d2732;
wire [40:0] d282,d284,d288,d2816,d2832;
wire [40:0] d292,d294,d298,d2916,d2932;
wire [40:0] d302,d304,d308,d3016,d3032;
wire [40:0] d312,d314,d318,d3116,d3132;

storage32_41 s00({o0s,o0},d002,d004,d008,d0016,d0032,se0,clk,reset);
storage32_41 s01({o1s,o1},d012,d014,d018,d0116,d0132,se1,clk,reset);
storage32_41 s02({o2s,o2},d022,d024,d028,d0216,d0232,se2,clk,reset);
storage32_41 s03({o3s,o3},d032,d034,d038,d0316,d0332,se3,clk,reset);
storage32_41 s04({o4s,o4},d042,d044,d048,d0416,d0432,se4,clk,reset);
storage32_41 s05({o5s,o5},d052,d054,d058,d0516,d0532,se5,clk,reset);
storage32_41 s06({o6s,o6},d062,d064,d068,d0616,d0632,se6,clk,reset);
storage32_41 s07({o7s,o7},d072,d074,d078,d0716,d0732,se7,clk,reset);
storage32_41 s08({o8s,o8},d082,d084,d088,d0816,d0832,se8,clk,reset);
storage32_41 s09({o9s,o9},d092,d094,d098,d0916,d0932,se9,clk,reset);
storage32_41 s10({o10s,o10},d102,d104,d108,d1016,d1032,se10,clk,reset);
storage32_41 s11({o11s,o11},d112,d114,d118,d1116,d1132,se11,clk,reset);
storage32_41 s12({o12s,o12},d122,d124,d128,d1216,d1232,se12,clk,reset);
storage32_41 s13({o13s,o13},d132,d134,d138,d1316,d1332,se13,clk,reset);
storage32_41 s14({o14s,o14},d142,d144,d148,d1416,d1432,se14,clk,reset);
storage32_41 s15({o15s,o15},d152,d154,d158,d1516,d1532,se15,clk,reset);
storage32_41 s16({o16s,o16},d162,d164,d168,d1616,d1632,se16,clk,reset);
storage32_41 s17({o17s,o17},d172,d174,d178,d1716,d1732,se17,clk,reset);
storage32_41 s18({o18s,o18},d182,d184,d188,d1816,d1832,se18,clk,reset);
storage32_41 s19({o19s,o19},d192,d194,d198,d1916,d1932,se19,clk,reset);
storage32_41 s20({o20s,o20},d202,d204,d208,d2016,d2032,se20,clk,reset);
storage32_41 s21({o21s,o21},d212,d214,d218,d2116,d2132,se21,clk,reset);
storage32_41 s22({o22s,o22},d222,d224,d228,d2216,d2232,se22,clk,reset);
storage32_41 s23({o23s,o23},d232,d234,d238,d2316,d2332,se23,clk,reset);
storage32_41 s24({o24s,o24},d242,d244,d248,d2416,d2432,se24,clk,reset);
storage32_41 s25({o25s,o25},d252,d254,d258,d2516,d2532,se25,clk,reset);
storage32_41 s26({o26s,o26},d262,d264,d268,d2616,d2632,se26,clk,reset);
storage32_41 s27({o27s,o27},d272,d274,d278,d2716,d2732,se27,clk,reset);
storage32_41 s28({o28s,o28},d282,d284,d288,d2816,d2832,se28,clk,reset);
storage32_41 s29({o29s,o29},d292,d294,d298,d2916,d2932,se29,clk,reset);
storage32_41 s30({o30s,o30},d302,d304,d308,d3016,d3032,se30,clk,reset);
storage32_41 s31({o31s,o31},d312,d314,d318,d3116,d3132,se31,clk,reset);

mux5_41 m00({oo0s,oo0},d002,d004,d008,d0016,d0032,se);
mux5_41 m01({oo1s,oo1},d012,d014,d018,d0116,d0132,se);
mux5_41 m02({oo2s,oo2},d022,d024,d028,d0216,d0232,se);
mux5_41 m03({oo3s,oo3},d032,d034,d038,d0316,d0332,se);
mux5_41 m04({oo4s,oo4},d042,d044,d048,d0416,d0432,se);
mux5_41 m05({oo5s,oo5},d052,d054,d058,d0516,d0532,se);
mux5_41 m06({oo6s,oo6},d062,d064,d068,d0616,d0632,se);
mux5_41 m07({oo7s,oo7},d072,d074,d078,d0716,d0732,se);
mux5_41 m08({oo8s,oo8},d082,d084,d088,d0816,d0832,se);
mux5_41 m09({oo9s,oo9},d092,d094,d098,d0916,d0932,se);
mux5_41 m10({oo10s,oo10},d102,d104,d108,d1016,d1032,se);
mux5_41 m11({oo11s,oo11},d112,d114,d118,d1116,d1132,se);
mux5_41 m12({oo12s,oo12},d122,d124,d128,d1216,d1232,se);
mux5_41 m13({oo13s,oo13},d132,d134,d138,d1316,d1332,se);
mux5_41 m14({oo14s,oo14},d142,d144,d148,d1416,d1432,se);
mux5_41 m15({oo15s,oo15},d152,d154,d158,d1516,d1532,se);
mux5_41 m16({oo16s,oo16},d162,d164,d168,d1616,d1632,se);
mux5_41 m17({oo17s,oo17},d172,d174,d178,d1716,d1732,se);
mux5_41 m18({oo18s,oo18},d182,d184,d188,d1816,d1832,se);
mux5_41 m19({oo19s,oo19},d192,d194,d198,d1916,d1932,se);
mux5_41 m20({oo20s,oo20},d202,d204,d208,d2016,d2032,se);
mux5_41 m21({oo21s,oo21},d212,d214,d218,d2116,d2132,se);
mux5_41 m22({oo22s,oo22},d222,d224,d228,d2216,d2232,se);
mux5_41 m23({oo23s,oo23},d232,d234,d238,d2316,d2332,se);
mux5_41 m24({oo24s,oo24},d242,d244,d248,d2416,d2432,se);
mux5_41 m25({oo25s,oo25},d252,d254,d258,d2516,d2532,se);
mux5_41 m26({oo26s,oo26},d262,d264,d268,d2616,d2632,se);
mux5_41 m27({oo27s,oo27},d272,d274,d278,d2716,d2732,se);
mux5_41 m28({oo28s,oo28},d282,d284,d288,d2816,d2832,se);
mux5_41 m29({oo29s,oo29},d292,d294,d298,d2916,d2932,se);
mux5_41 m30({oo30s,oo30},d302,d304,d308,d3016,d3032,se);
mux5_41 m31({oo31s,oo31},d312,d314,d318,d3116,d3132,se);

endmodule


//32 number of 5-to-1 multiplexers used for input of 32x32 buffer in proposed Interger DCT folded architecture

//`include "mux5to1_41.v"

module col_mux_inp_buf_folded_pro(

ou20s,ou21s,ou22s,ou23s,ou24s,ou25s,ou26s,ou27s,ou28s,ou29s,ou210s,ou211s,ou212s,ou213s,ou214s,ou215s,
ou40s,ou41s,ou42s,ou43s,ou44s,ou45s,ou46s,ou47s,
ou80s,ou81s,ou82s,ou83s,
ou160s,ou161s,
ou320s,

ou20,ou21,ou22,ou23,ou24,ou25,ou26,ou27,ou28,ou29,ou210,ou211,ou212,ou213,ou214,ou215,
ou40,ou41,ou42,ou43,ou44,ou45,ou46,ou47,
ou80,ou81,ou82,ou83,
ou160,ou161,
ou320,

se,

o0s,o1s,o2s,o3s,o4s,o5s,o6s,o7s,o8s,o9s,o10s,o11s,o12s,o13s,o14s,o15s,o16s,o17s,o18s,o19s,o20s,o21s,o22s,o23s,o24s,o25s,o26s,o27s,o28s,o29s,o30s,o31s,
o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,o10,o11,o12,o13,o14,o15,o16,o17,o18,o19,o20,o21,o22,o23,o24,o25,o26,o27,o28,o29,o30,o31

);

input ou20s,ou21s,ou22s,ou23s,ou24s,ou25s,ou26s,ou27s,ou28s,ou29s,ou210s,ou211s,ou212s,ou213s,ou214s,ou215s,
ou40s,ou41s,ou42s,ou43s,ou44s,ou45s,ou46s,ou47s,
ou80s,ou81s,ou82s,ou83s,
ou160s,ou161s,
ou320s;

input [39:0] ou20,ou21,ou22,ou23,ou24,ou25,ou26,ou27,ou28,ou29,ou210,ou211,ou212,ou213,ou214,ou215,
ou40,ou41,ou42,ou43,ou44,ou45,ou46,ou47,
ou80,ou81,ou82,ou83,
ou160,ou161,
ou320;

input [2:0] se;

output [39:0] o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,o10,o11,o12,o13,o14,o15,o16,o17,o18,o19,o20,o21,o22,o23,o24,o25,o26,o27,o28,o29,o30,o31;
output o0s,o1s,o2s,o3s,o4s,o5s,o6s,o7s,o8s,o9s,o10s,o11s,o12s,o13s,o14s,o15s,o16s,o17s,o18s,o19s,o20s,o21s,o22s,o23s,o24s,o25s,o26s,o27s,o28s,o29s,o30s,o31s;

mux5to1_41 m00({o0s,o0},{ou320s,ou320},{ou160s,ou160},{ou80s,ou80},{ou40s,ou40},{ou20s,ou20},se);
mux5to1_41 m01({o1s,o1},{ou320s,ou320},{ou160s,ou160},{ou80s,ou80},{ou40s,ou40},{ou20s,ou20},se);
mux5to1_41 m02({o2s,o2},{ou320s,ou320},{ou160s,ou160},{ou80s,ou80},{ou40s,ou40},{ou21s,ou21},se);
mux5to1_41 m03({o3s,o3},{ou320s,ou320},{ou160s,ou160},{ou80s,ou80},{ou40s,ou40},{ou21s,ou21},se);
mux5to1_41 m04({o4s,o4},{ou320s,ou320},{ou160s,ou160},{ou80s,ou80},{ou41s,ou41},{ou22s,ou22},se);
mux5to1_41 m05({o5s,o5},{ou320s,ou320},{ou160s,ou160},{ou80s,ou80},{ou41s,ou41},{ou22s,ou22},se);
mux5to1_41 m06({o6s,o6},{ou320s,ou320},{ou160s,ou160},{ou80s,ou80},{ou41s,ou41},{ou23s,ou23},se);
mux5to1_41 m07({o7s,o7},{ou320s,ou320},{ou160s,ou160},{ou80s,ou80},{ou41s,ou41},{ou23s,ou23},se);
mux5to1_41 m08({o8s,o8},{ou320s,ou320},{ou160s,ou160},{ou81s,ou81},{ou42s,ou42},{ou24s,ou24},se);
mux5to1_41 m09({o9s,o9},{ou320s,ou320},{ou160s,ou160},{ou81s,ou81},{ou42s,ou42},{ou24s,ou24},se);
mux5to1_41 m010({o10s,o10},{ou320s,ou320},{ou160s,ou160},{ou81s,ou81},{ou42s,ou42},{ou25s,ou25},se);
mux5to1_41 m011({o11s,o11},{ou320s,ou320},{ou160s,ou160},{ou81s,ou81},{ou42s,ou42},{ou25s,ou25},se);
mux5to1_41 m012({o12s,o12},{ou320s,ou320},{ou160s,ou160},{ou81s,ou81},{ou43s,ou43},{ou26s,ou26},se);
mux5to1_41 m013({o13s,o13},{ou320s,ou320},{ou160s,ou160},{ou81s,ou81},{ou43s,ou43},{ou26s,ou26},se);
mux5to1_41 m014({o14s,o14},{ou320s,ou320},{ou160s,ou160},{ou81s,ou81},{ou43s,ou43},{ou27s,ou27},se);
mux5to1_41 m015({o15s,o15},{ou320s,ou320},{ou160s,ou160},{ou81s,ou81},{ou43s,ou43},{ou27s,ou27},se);
mux5to1_41 m016({o16s,o16},{ou320s,ou320},{ou161s,ou161},{ou82s,ou82},{ou44s,ou44},{ou28s,ou28},se);
mux5to1_41 m017({o17s,o17},{ou320s,ou320},{ou161s,ou161},{ou82s,ou82},{ou44s,ou44},{ou28s,ou28},se);
mux5to1_41 m018({o18s,o18},{ou320s,ou320},{ou161s,ou161},{ou82s,ou82},{ou44s,ou44},{ou29s,ou29},se);
mux5to1_41 m019({o19s,o19},{ou320s,ou320},{ou161s,ou161},{ou82s,ou82},{ou44s,ou44},{ou29s,ou29},se);
mux5to1_41 m020({o20s,o20},{ou320s,ou320},{ou161s,ou161},{ou82s,ou82},{ou45s,ou45},{ou210s,ou210},se);
mux5to1_41 m021({o21s,o21},{ou320s,ou320},{ou161s,ou161},{ou82s,ou82},{ou45s,ou45},{ou210s,ou210},se);
mux5to1_41 m022({o22s,o22},{ou320s,ou320},{ou161s,ou161},{ou82s,ou82},{ou45s,ou45},{ou211s,ou211},se);
mux5to1_41 m023({o23s,o23},{ou320s,ou320},{ou161s,ou161},{ou82s,ou82},{ou45s,ou45},{ou211s,ou211},se);
mux5to1_41 m024({o24s,o24},{ou320s,ou320},{ou161s,ou161},{ou83s,ou83},{ou46s,ou46},{ou212s,ou212},se);
mux5to1_41 m025({o25s,o25},{ou320s,ou320},{ou161s,ou161},{ou83s,ou83},{ou46s,ou46},{ou212s,ou212},se);
mux5to1_41 m026({o26s,o26},{ou320s,ou320},{ou161s,ou161},{ou83s,ou83},{ou46s,ou46},{ou213s,ou213},se);
mux5to1_41 m027({o27s,o27},{ou320s,ou320},{ou161s,ou161},{ou83s,ou83},{ou46s,ou46},{ou213s,ou213},se);
mux5to1_41 m028({o28s,o28},{ou320s,ou320},{ou161s,ou161},{ou83s,ou83},{ou47s,ou47},{ou214s,ou214},se);
mux5to1_41 m029({o29s,o29},{ou320s,ou320},{ou161s,ou161},{ou83s,ou83},{ou47s,ou47},{ou214s,ou214},se);
mux5to1_41 m030({o30s,o30},{ou320s,ou320},{ou161s,ou161},{ou83s,ou83},{ou47s,ou47},{ou215s,ou215},se);
mux5to1_41 m031({o31s,o31},{ou320s,ou320},{ou161s,ou161},{ou83s,ou83},{ou47s,ou47},{ou215s,ou215},se);

endmodule


//mux5 to 1

module mux5to1_41(o,o1,o2,o3,o4,o5,dir);

input [2:0] dir;
input [40:0] o1,o2,o3,o4,o5;
output [40:0] o;

reg [40:0] o;

always@(o1 or o2 or o3 or o4 or o5 or dir)
	begin
	 case(dir)
	  3'b000: o=o1;
	  3'b001: o=o2;
	  3'b010: o=o3;
	  3'b011: o=o4;
	  3'b100: o=o5;	  
	default: o = 1'bx;
	 endcase
	end

endmodule



// storage buffer

//`include "mux2to1_41.v"
//`include "dflipflop41.v"

module storage32_41(i,d32,s,clk,reset);

input [40:0] i;
input s,clk,reset;//s is 0 for feed back and 1 for feed forward
output [40:0] d32;

wire [40:0] m1,m2,m3,m4,m5,m6,m7,m8,m9,m10,m11,m12,m13,m14,m15,m16,m17,m18,m19,m20,m21,m22,m23,m24,m25,m26,m27,m28,m29,m30,m31,m32;
wire [40:0] d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28,d29,d30,d31,d32;

mux2to1_41 mu1(m1,d1,i,s); 
dflipflop41 df1(d1,m1,clk,reset);

mux2to1_41 mu2(m2,d2,d1,s);
dflipflop41 df2(d2,m2,clk,reset);

mux2to1_41 mu3(m3,d3,d2,s);
dflipflop41 df3(d3,m3,clk,reset);

mux2to1_41 mu4(m4,d4,d3,s);
dflipflop41 df4(d4,m4,clk,reset);

mux2to1_41 mu5(m5,d5,d4,s);
dflipflop41 df5(d5,m5,clk,reset);

mux2to1_41 mu6(m6,d6,d5,s);
dflipflop41 df6(d6,m6,clk,reset);

mux2to1_41 mu7(m7,d7,d6,s);
dflipflop41 df7(d7,m7,clk,reset);

mux2to1_41 mu8(m8,d8,d7,s);
dflipflop41 df8(d8,m8,clk,reset);

mux2to1_41 mu9(m9,d9,d8,s);
dflipflop41 df9(d9,m9,clk,reset);

mux2to1_41 mu10(m10,d10,d9,s);
dflipflop41 df10(d10,m10,clk,reset);

mux2to1_41 mu11(m11,d11,d10,s);
dflipflop41 df11(d11,m11,clk,reset);

mux2to1_41 mu12(m12,d12,d11,s);
dflipflop41 df12(d12,m12,clk,reset);

mux2to1_41 mu13(m13,d13,d12,s);
dflipflop41 df13(d13,m13,clk,reset);

mux2to1_41 mu14(m14,d14,d13,s);
dflipflop41 df14(d14,m14,clk,reset);

mux2to1_41 mu15(m15,d15,d14,s);
dflipflop41 df15(d15,m15,clk,reset);

mux2to1_41 mu16(m16,d16,d15,s);
dflipflop41 df16(d16,m16,clk,reset);

mux2to1_41 mu17(m17,d17,d16,s);
dflipflop41 df17(d17,m17,clk,reset);

mux2to1_41 mu18(m18,d18,d17,s);
dflipflop41 df18(d18,m18,clk,reset);

mux2to1_41 mu19(m19,d19,d18,s);
dflipflop41 df19(d19,m19,clk,reset);

mux2to1_41 mu20(m20,d20,d19,s);
dflipflop41 df20(d20,m20,clk,reset);

mux2to1_41 mu21(m21,d21,d20,s);
dflipflop41 df21(d21,m21,clk,reset);

mux2to1_41 mu22(m22,d22,d21,s);
dflipflop41 df22(d22,m22,clk,reset);

mux2to1_41 mu23(m23,d23,d22,s);
dflipflop41 df23(d23,m23,clk,reset);

mux2to1_41 mu24(m24,d24,d23,s);
dflipflop41 df24(d24,m24,clk,reset);

mux2to1_41 mu25(m25,d25,d24,s);
dflipflop41 df25(d25,m25,clk,reset);

mux2to1_41 mu26(m26,d26,d25,s);
dflipflop41 df26(d26,m26,clk,reset);

mux2to1_41 mu27(m27,d27,d26,s);
dflipflop41 df27(d27,m27,clk,reset);

mux2to1_41 mu28(m28,d28,d27,s);
dflipflop41 df28(d28,m28,clk,reset);

mux2to1_41 mu29(m29,d29,d28,s);
dflipflop41 df29(d29,m29,clk,reset);

mux2to1_41 mu30(m30,d30,d29,s);
dflipflop41 df30(d30,m30,clk,reset);

mux2to1_41 mu31(m31,d31,d30,s);
dflipflop41 df31(d31,m31,clk,reset);

mux2to1_41 mu32(m32,d32,d31,s);
dflipflop41 df32(d32,m32,clk,reset);

endmodule

//mux5 to 1

module mux5_41(o,o1,o2,o3,o4,o5,dir);

input [2:0] dir;
input [40:0] o1,o2,o3,o4,o5;
output [40:0] o;

reg [40:0] o;

always@(o1 or o2 or o3 or o4 or o5 or dir)
	begin
	 case(dir)
	  3'b000: o=o5;
	  3'b001: o=o4;
	  3'b010: o=o3;
	  3'b011: o=o2;
	  3'b100: o=o1;	  
	default: o = 25'bx;
	 endcase
	end

endmodule

//2 to 1 multiplexer design

module mux2to1_41(out,i1,i2,s);

input [40:0] i1,i2;
input s;
output [40:0] out;
reg [40:0] out;

always@(i1 or i2 or s)
	begin
	 case(s)
	  1'b0:out=i1;
	  1'b1:out=i2;
	 endcase
	end

endmodule

// D flip flop

module dflipflop41(q,d,clk,reset);
output [40:0] q;
input [40:0] d;
input clk,reset;
reg [40:0] q;
always@(posedge reset or negedge clk)
if(reset)
q<=41'b00000000;
else
q<=d;
endmodule




















`default_nettype wire
